module hello2;
  initial
    begin
      $display("Hello, World 2");
      $finish ;
    end
endmodule
