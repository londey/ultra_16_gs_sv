

module top (
    // Add your module ports here
);
     
// Add your module implementation here
     
endmodule
    port_list
);
